`timescale 1 ns / 1 ps

module mdunit(input         clk, reset,
              input  [31:0] srca, srcb,
              input  [2:0]  alushcontrol,
              input         mdstart, 
              output [31:0] data_out,
              output        mdrun);
    
endmodule

